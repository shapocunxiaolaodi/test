module design1(
	input clk,
	output clk_3div
);

endmodule;
