module design1(
);

endmodule;
