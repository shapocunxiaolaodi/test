module design1(
  input clk
);

endmodule;
